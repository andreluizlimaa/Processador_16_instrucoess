library verilog;
use verilog.vl_types.all;
entity Comparator_LG_1bit_vlg_check_tst is
    port(
        e               : in     vl_logic;
        g               : in     vl_logic;
        l               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Comparator_LG_1bit_vlg_check_tst;
