library verilog;
use verilog.vl_types.all;
entity Right_Shifter_vlg_vec_tst is
end Right_Shifter_vlg_vec_tst;
