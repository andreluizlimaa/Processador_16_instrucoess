library verilog;
use verilog.vl_types.all;
entity Mux4x1_16bit_vlg_vec_tst is
end Mux4x1_16bit_vlg_vec_tst;
