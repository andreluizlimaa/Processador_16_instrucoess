library verilog;
use verilog.vl_types.all;
entity Adder_16bit_vlg_vec_tst is
end Adder_16bit_vlg_vec_tst;
