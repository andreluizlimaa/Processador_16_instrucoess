library verilog;
use verilog.vl_types.all;
entity Mux2x1_16bit_vlg_vec_tst is
end Mux2x1_16bit_vlg_vec_tst;
