library verilog;
use verilog.vl_types.all;
entity Comparator_LG_16bit_vlg_check_tst is
    port(
        G               : in     vl_logic;
        L               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Comparator_LG_16bit_vlg_check_tst;
