library verilog;
use verilog.vl_types.all;
entity Comparator_LG_1bit_vlg_vec_tst is
end Comparator_LG_1bit_vlg_vec_tst;
