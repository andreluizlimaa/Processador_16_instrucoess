library verilog;
use verilog.vl_types.all;
entity Left_Shifter_vlg_vec_tst is
end Left_Shifter_vlg_vec_tst;
