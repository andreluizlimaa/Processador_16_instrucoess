library verilog;
use verilog.vl_types.all;
entity flipflopD2_vlg_vec_tst is
end flipflopD2_vlg_vec_tst;
