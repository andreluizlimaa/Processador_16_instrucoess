library ieee;
use ieee.std_logic_1164.all;

ENTITY Decode_4x16 IS
PORT(
    A3, A2, A1, A0, E: IN std_logic;
    Y15, Y14, Y13, Y12, Y11, Y10, Y9, Y8, Y7, Y6, Y5, Y4, Y3, Y2, Y1, Y0 : OUT std_logic
);
END ENTITY;

ARCHITECTURE comb OF Decode_4x16 IS
BEGIN
    Y0 <= E AND NOT(A3) AND NOT(A2) AND NOT(A1) AND NOT(A0);
    Y1 <= E AND NOT(A3) AND NOT(A2) AND NOT(A1) AND A0;
    Y2 <= E AND NOT(A3) AND NOT(A2) AND A1 AND NOT(A0);
    Y3 <= E AND NOT(A3) AND NOT(A2) AND A1 AND A0;
    Y4 <= E AND NOT(A3) AND A2 AND NOT(A1) AND NOT(A0);
    Y5 <= E AND NOT(A3) AND A2 AND NOT(A1) AND A0;
    Y6 <= E AND NOT(A3) AND A2 AND A1 AND NOT(A0);
    Y7 <= E AND NOT(A3) AND A2 AND A1 AND A0;
    Y8 <= E AND A3 AND NOT(A2) AND NOT(A1) AND NOT(A0);
    Y9 <= E AND A3 AND NOT(A2) AND NOT(A1) AND A0;
    Y10 <= E AND A3 AND NOT(A2) AND A1 AND NOT(A0);
    Y11 <= E AND A3 AND NOT(A2) AND A1 AND A0;
    Y12 <= E AND A3 AND A2 AND NOT(A1) AND NOT(A0);
    Y13 <= E AND A3 AND A2 AND NOT(A1) AND A0;
    Y14 <= E AND A3 AND A2 AND A1 AND NOT(A0);
    Y15 <= E AND A3 AND A2 AND A1 AND A0;
END ARCHITECTURE;
