library verilog;
use verilog.vl_types.all;
entity Mux16x1_1bit_vlg_vec_tst is
end Mux16x1_1bit_vlg_vec_tst;
