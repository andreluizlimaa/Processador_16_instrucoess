library verilog;
use verilog.vl_types.all;
entity Inst_Reg_vlg_vec_tst is
end Inst_Reg_vlg_vec_tst;
