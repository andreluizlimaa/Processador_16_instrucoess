library verilog;
use verilog.vl_types.all;
entity Program_Counter_vlg_vec_tst is
end Program_Counter_vlg_vec_tst;
