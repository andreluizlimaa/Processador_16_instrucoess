library verilog;
use verilog.vl_types.all;
entity FlipFlopD2_vlg_vec_tst is
end FlipFlopD2_vlg_vec_tst;
