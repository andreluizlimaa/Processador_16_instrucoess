library verilog;
use verilog.vl_types.all;
entity FlipflopD_vlg_vec_tst is
end FlipflopD_vlg_vec_tst;
