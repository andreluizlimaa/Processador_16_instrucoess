library verilog;
use verilog.vl_types.all;
entity Mux16x1_1bit_vlg_check_tst is
    port(
        O               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Mux16x1_1bit_vlg_check_tst;
